`timescale 1us/1us

module round_robin_arbiter (
  input     logic          clk  ,
  input     logic          reset,

  input     logic   [3:0]  req_i,
  output    logic   [3:0]  gnt_o
);

//insert the logic here

endmodule